----------
-- File Name : Pattern_8_slv.vhd
-- Function : Display the Input Pattern on the 7 Segment LED
-- Author : Manabu Inoue
-- Rev and Date : 1.0 , 2008/10/19 , original source
----------


library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_signed.all;


entity Pattern_8_slv is

	port (
		SW : in std_logic_vector(2 downto 0);
		SEG7 : out std_logic_vector(6 downto 0)
	);

end Pattern_8_slv;


architecture RTL of Pattern_8_slv is





begin





end RTL;